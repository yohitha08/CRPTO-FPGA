module expansion(input[1:32] right,output[0:47] exp);
assign exp[0]=right[32];
assign exp[1]=right[1];
assign exp[2]=right[2];
assign exp[3]=right[3];
assign exp[4]=right[4];
assign exp[5]=right[5];
assign exp[6]=right[4];
assign exp[7]=right[5];
assign exp[8]=right[6];
assign exp[9]=right[7];
assign exp[10]=right[8];
assign exp[11]=right[9];
assign exp[12]=right[8];
assign exp[13]=right[9];
assign exp[14]=right[10];
assign exp[15]=right[11];
assign exp[16]=right[12];
assign exp[17]=right[13];
assign exp[18]=right[12];
assign exp[19]=right[13];
assign exp[20]=right[14];
assign exp[21]=right[15];
assign exp[22]=right[16];
assign exp[23]=right[17];
assign exp[24]=right[16];
assign exp[25]=right[17];
assign exp[26]=right[18];
assign exp[27]=right[19];
assign exp[28]=right[20];
assign exp[29]=right[21];
assign exp[30]=right[20];
assign exp[31]=right[21];
assign exp[32]=right[22];
assign exp[33]=right[23];
assign exp[34]=right[24];
assign exp[35]=right[25];
assign exp[36]=right[24];
assign exp[37]=right[25];
assign exp[38]=right[26];
assign exp[39]=right[27];
assign exp[40]=right[28];
assign exp[41]=right[29];
assign exp[42]=right[28];
assign exp[43]=right[29];
assign exp[44]=right[30];
assign exp[45]=right[31];
assign exp[46]=right[32];
assign exp[47]=right[1];
endmodule
